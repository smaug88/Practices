--
-- DLX_PROG2.vhd
--
-- Programa para el DLX32p
-- Se ha insertado nop para evitar las dependencias. Esta es la diferencia con DLX_PROG.vhd
-- que es el que se ha utilizado para DLX32s monociclo.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
use work.DLX_pack.all;

package DLX_prog2 is
  type ROM_TABLE is array (0 to 29) of ROM_WORD;

  constant ROM: ROM_TABLE := ROM_TABLE'(

      ROM_WORD'("00110100000111100000000000000000"),
      ROM_WORD'("00110100000010110000000000000001"),
      ROM_WORD'("00110100000000010000000000000110"),
      ROM_WORD'("00110100000000100000000000001011"),
      ROM_WORD'("00110100000000110000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000010010110010000000100100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000100000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000010001100000100000"),
      ROM_WORD'("00000000010010110001000000000111"),
      ROM_WORD'("00000000001010110000100000000100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000010000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000000001100000100000")
      );

end DLX_prog2;
