--
-- DLX_PROG2.vhd
--
-- Programa para el DLX32p
-- Se ha insertado nop para evitar las dependencias. Esta es la diferencia con DLX_PROG.vhd
-- que es el que se ha utilizado para DLX32s monociclo.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
use work.DLX_pack.all;

package DLX_prog2 is
  type ROM_TABLE is array (0 to 170) of ROM_WORD;

  constant ROM: ROM_TABLE := ROM_TABLE'(

      ROM_WORD'("00110100000111100000000000000000"),
      ROM_WORD'("00110100000000110000000000000000"),
      ROM_WORD'("00110100000010100001111100100000"),
      ROM_WORD'("00110100000011000000011100100000"),
      ROM_WORD'("00110100000010110000000000000001"),
      ROM_WORD'("00110100000011100000000011111111"),
      ROM_WORD'("00110100000011010000000000001000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000001010011100000100000100100"),
      ROM_WORD'("00000001100011100001000000100100"),
      ROM_WORD'("00001000000000000000000000100000"),
      ROM_WORD'("00000001010011010101000000000111"),
      ROM_WORD'("00000001100011010110000000000111"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010001010000000000000001011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000010010110010000000100100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000100000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000010001100000100000"),
      ROM_WORD'("00000000010010110001000000000111"),
      ROM_WORD'("00000000001010110000100000000100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000010000001111111110101100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00110100000010100010000100100000"),
      ROM_WORD'("00110100000011000000110100001000"),
      ROM_WORD'("00110100000010110000000000000001"),
      ROM_WORD'("00000001010011100000100000100100"),
      ROM_WORD'("00000001100011100001000000100100"),
      ROM_WORD'("00001000000000000000000000100000"),
      ROM_WORD'("00000001010011010101000000000111"),
      ROM_WORD'("00000001100011010110000000000111"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010001010000000000000001011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000010010110010000000100100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000100000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000010001100000100000"),
      ROM_WORD'("00000000010010110001000000000111"),
      ROM_WORD'("00000000001010110000100000000100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000010000001111111110101100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00110100000010100001111100100000"),
      ROM_WORD'("00110100000011000001100100101100"),
      ROM_WORD'("00110100000010110000000000000001"),
      ROM_WORD'("00000001010011100000100000100100"),
      ROM_WORD'("00000001100011100001000000100100"),
      ROM_WORD'("00001000000000000000000000100000"),
      ROM_WORD'("00000001010011010101000000000111"),
      ROM_WORD'("00000001100011010110000000000111"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010001010000000000000001011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000010010110010000000100100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000100000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000010001100000100000"),
      ROM_WORD'("00000000010010110001000000000111"),
      ROM_WORD'("00000000001010110000100000000100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000010000001111111110101100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00110100000010100010000100100000"),
      ROM_WORD'("00110100000011000000001000001011"),
      ROM_WORD'("00110100000010110000000000000001"),
      ROM_WORD'("00000001010011100000100000100100"),
      ROM_WORD'("00000001100011100001000000100100"),
      ROM_WORD'("00001000000000000000000000100000"),
      ROM_WORD'("00000001010011010101000000000111"),
      ROM_WORD'("00000001100011010110000000000111"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010001010000000000000001011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000010010110010000000100100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000100000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000010001100000100000"),
      ROM_WORD'("00000000010010110001000000000111"),
      ROM_WORD'("00000000001010110000100000000100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000010000001111111110101100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00110100000010100001111100100000"),
      ROM_WORD'("00110100000011000000100100010001"),
      ROM_WORD'("00110100000010110000000000000001"),
      ROM_WORD'("00000001010011100000100000100100"),
      ROM_WORD'("00000001100011100001000000100100"),
      ROM_WORD'("00001000000000000000000000100000"),
      ROM_WORD'("00000001010011010101000000000111"),
      ROM_WORD'("00000001100011010110000000000111"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010001010000000000000001011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111011000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000010010110010000000100100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000100000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011000010001100000100000"),
      ROM_WORD'("00000000010010110001000000000111"),
      ROM_WORD'("00000000001010110000100000000100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00010000010000001111111110101100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000")
      );

end DLX_prog2;
