--
-- DLX_PROG2.vhd
--
-- Programa para el DLX32p
-- Se ha insertado nop para evitar las dependencias. Esta es la diferencia con DLX_PROG.vhd
-- que es el que se ha utilizado para DLX32s monociclo.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
use work.DLX_pack.all;

package DLX_prog2 is
  type ROM_TABLE is array (0 to 40) of ROM_WORD;

  constant ROM: ROM_TABLE := ROM_TABLE'(

      ROM_WORD'("00110100000111100000000000000000"),
      ROM_WORD'("00110100000000010000000000001010"),
      ROM_WORD'("00001100000000000000000000001100"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00001011111111111111111111110000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("10101111110000100000000000000000"),
      ROM_WORD'("00110100000000100000000000000001"),
      ROM_WORD'("00000011110000101111000000100000"),
      ROM_WORD'("10101111110000010000000000000000"),
      ROM_WORD'("00000011110000101111000000100000"),
      ROM_WORD'("10101111110000110000000000000000"),
      ROM_WORD'("00000011110000101111000000100000"),
      ROM_WORD'("10101111110111110000000000000000"),
      ROM_WORD'("00000011110000101111000000100000"),
      ROM_WORD'("00110100000000100000000000000010"),
      ROM_WORD'("00000000001000100001000000101010"),
      ROM_WORD'("00010000010000000000000000001100"),
      ROM_WORD'("00000000000000010101100000100000"),
      ROM_WORD'("00001000000000000000000000101000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00110100000000100000000000000001"),
      ROM_WORD'("00000000001000100000100000100010"),
      ROM_WORD'("00001111111111111111111110111000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000000010110001100000100000"),
      ROM_WORD'("00000000001000100000100000100010"),
      ROM_WORD'("00001111111111111111111110101000"),
      ROM_WORD'("00000000000000000000000000000000"),
      ROM_WORD'("00000000011010110101100000100000"),
      ROM_WORD'("00110100000000100000000000000001"),
      ROM_WORD'("00000011110000101111000000100010"),
      ROM_WORD'("10001111110111110000000000000000"),
      ROM_WORD'("00000011110000101111000000100010"),
      ROM_WORD'("10001111110000110000000000000000"),
      ROM_WORD'("00000011110000101111000000100010"),
      ROM_WORD'("10001111110000010000000000000000"),
      ROM_WORD'("00000011110000101111000000100010"),
      ROM_WORD'("10001111110000100000000000000000"),
      ROM_WORD'("01001011111000000000000000000000"),
      ROM_WORD'("00000000000000000000000000000000")
      );

end DLX_prog2;
